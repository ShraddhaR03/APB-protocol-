package apb_pkg;
`include "uvm_macros.svh" 
import uvm_pkg::*;

`include "seq_item.sv"
`include "slave_monitor.sv"
`include "master_monitor.sv"
`include "apb_driver.sv"
`include "master_seqr.sv"
`include "master_agent_config.sv"
`include "slave_agent_config.sv"
`include "env_config.sv"
`include "slave_agent.sv"
`include "master_agent.sv"
`include "scoreboard.sv"
`include "coverage_collector.sv"

`include "apb_vseqr.sv"
`include "apb_env.sv"
 `include "apb_seq.sv"
`include "apb_vseq.sv"
 `include "apb_test.sv"

endpackage